`include "types.vh"


module alu (


    
);

endmodule