import testbench_pkg::*;

class interface_tester extends base_testbench;

    task tb_setup();
        super.tb_setup();
    endtask

    virtual task run();
        super.run();
    endtask 


endclass