module core (
    input  clk,    // Clock
    input  rst_n,  // Asynchronous reset active low
    input  i_data,
    output i_addr,
    input  d_data,
    output d_addr,
    output o_data,
    output wr_en,
    output rd_en
);

endmodule