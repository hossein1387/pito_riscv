`include "types.svh"
`include "instr.svh"
