`include "types.svh"
`include "instr.svh"

module decoder (
    input clk,    // Clock
    input i_data, // Clock Enable
    i
);

endmodule