../utils/utils.sv